    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   SaveData   	positionX	positionY	positionZcurrentSceneIDnamedataTime        ��B    33EB      Alexsmithcore�fx�ֈ